// HPS.v

// Generated using ACDS version 17.0 595

`timescale 1 ps / 1 ps
module HPS (
		input  wire        clk_clk,                                          //                    clk.clk
		input  wire        hps_f2h_axi_clock_clk,                            //      hps_f2h_axi_clock.clk
		input  wire [7:0]  hps_f2h_axi_slave_awid,                           //      hps_f2h_axi_slave.awid
		input  wire [31:0] hps_f2h_axi_slave_awaddr,                         //                       .awaddr
		input  wire [3:0]  hps_f2h_axi_slave_awlen,                          //                       .awlen
		input  wire [2:0]  hps_f2h_axi_slave_awsize,                         //                       .awsize
		input  wire [1:0]  hps_f2h_axi_slave_awburst,                        //                       .awburst
		input  wire [1:0]  hps_f2h_axi_slave_awlock,                         //                       .awlock
		input  wire [3:0]  hps_f2h_axi_slave_awcache,                        //                       .awcache
		input  wire [2:0]  hps_f2h_axi_slave_awprot,                         //                       .awprot
		input  wire        hps_f2h_axi_slave_awvalid,                        //                       .awvalid
		output wire        hps_f2h_axi_slave_awready,                        //                       .awready
		input  wire [4:0]  hps_f2h_axi_slave_awuser,                         //                       .awuser
		input  wire [7:0]  hps_f2h_axi_slave_wid,                            //                       .wid
		input  wire [31:0] hps_f2h_axi_slave_wdata,                          //                       .wdata
		input  wire [3:0]  hps_f2h_axi_slave_wstrb,                          //                       .wstrb
		input  wire        hps_f2h_axi_slave_wlast,                          //                       .wlast
		input  wire        hps_f2h_axi_slave_wvalid,                         //                       .wvalid
		output wire        hps_f2h_axi_slave_wready,                         //                       .wready
		output wire [7:0]  hps_f2h_axi_slave_bid,                            //                       .bid
		output wire [1:0]  hps_f2h_axi_slave_bresp,                          //                       .bresp
		output wire        hps_f2h_axi_slave_bvalid,                         //                       .bvalid
		input  wire        hps_f2h_axi_slave_bready,                         //                       .bready
		input  wire [7:0]  hps_f2h_axi_slave_arid,                           //                       .arid
		input  wire [31:0] hps_f2h_axi_slave_araddr,                         //                       .araddr
		input  wire [3:0]  hps_f2h_axi_slave_arlen,                          //                       .arlen
		input  wire [2:0]  hps_f2h_axi_slave_arsize,                         //                       .arsize
		input  wire [1:0]  hps_f2h_axi_slave_arburst,                        //                       .arburst
		input  wire [1:0]  hps_f2h_axi_slave_arlock,                         //                       .arlock
		input  wire [3:0]  hps_f2h_axi_slave_arcache,                        //                       .arcache
		input  wire [2:0]  hps_f2h_axi_slave_arprot,                         //                       .arprot
		input  wire        hps_f2h_axi_slave_arvalid,                        //                       .arvalid
		output wire        hps_f2h_axi_slave_arready,                        //                       .arready
		input  wire [4:0]  hps_f2h_axi_slave_aruser,                         //                       .aruser
		output wire [7:0]  hps_f2h_axi_slave_rid,                            //                       .rid
		output wire [31:0] hps_f2h_axi_slave_rdata,                          //                       .rdata
		output wire [1:0]  hps_f2h_axi_slave_rresp,                          //                       .rresp
		output wire        hps_f2h_axi_slave_rlast,                          //                       .rlast
		output wire        hps_f2h_axi_slave_rvalid,                         //                       .rvalid
		input  wire        hps_f2h_axi_slave_rready,                         //                       .rready
		input  wire        hps_f2h_boot_from_fpga_boot_from_fpga_ready,      // hps_f2h_boot_from_fpga.boot_from_fpga_ready
		input  wire        hps_f2h_boot_from_fpga_boot_from_fpga_on_failure, //                       .boot_from_fpga_on_failure
		output wire        hps_h2f_reset_reset_n,                            //          hps_h2f_reset.reset_n
		output wire        hps_io_hps_io_emac1_inst_TX_CLK,                  //                 hps_io.hps_io_emac1_inst_TX_CLK
		output wire        hps_io_hps_io_emac1_inst_TXD0,                    //                       .hps_io_emac1_inst_TXD0
		output wire        hps_io_hps_io_emac1_inst_TXD1,                    //                       .hps_io_emac1_inst_TXD1
		output wire        hps_io_hps_io_emac1_inst_TXD2,                    //                       .hps_io_emac1_inst_TXD2
		output wire        hps_io_hps_io_emac1_inst_TXD3,                    //                       .hps_io_emac1_inst_TXD3
		input  wire        hps_io_hps_io_emac1_inst_RXD0,                    //                       .hps_io_emac1_inst_RXD0
		inout  wire        hps_io_hps_io_emac1_inst_MDIO,                    //                       .hps_io_emac1_inst_MDIO
		output wire        hps_io_hps_io_emac1_inst_MDC,                     //                       .hps_io_emac1_inst_MDC
		input  wire        hps_io_hps_io_emac1_inst_RX_CTL,                  //                       .hps_io_emac1_inst_RX_CTL
		output wire        hps_io_hps_io_emac1_inst_TX_CTL,                  //                       .hps_io_emac1_inst_TX_CTL
		input  wire        hps_io_hps_io_emac1_inst_RX_CLK,                  //                       .hps_io_emac1_inst_RX_CLK
		input  wire        hps_io_hps_io_emac1_inst_RXD1,                    //                       .hps_io_emac1_inst_RXD1
		input  wire        hps_io_hps_io_emac1_inst_RXD2,                    //                       .hps_io_emac1_inst_RXD2
		input  wire        hps_io_hps_io_emac1_inst_RXD3,                    //                       .hps_io_emac1_inst_RXD3
		inout  wire        hps_io_hps_io_sdio_inst_CMD,                      //                       .hps_io_sdio_inst_CMD
		inout  wire        hps_io_hps_io_sdio_inst_D0,                       //                       .hps_io_sdio_inst_D0
		inout  wire        hps_io_hps_io_sdio_inst_D1,                       //                       .hps_io_sdio_inst_D1
		output wire        hps_io_hps_io_sdio_inst_CLK,                      //                       .hps_io_sdio_inst_CLK
		inout  wire        hps_io_hps_io_sdio_inst_D2,                       //                       .hps_io_sdio_inst_D2
		inout  wire        hps_io_hps_io_sdio_inst_D3,                       //                       .hps_io_sdio_inst_D3
		inout  wire        hps_io_hps_io_usb1_inst_D0,                       //                       .hps_io_usb1_inst_D0
		inout  wire        hps_io_hps_io_usb1_inst_D1,                       //                       .hps_io_usb1_inst_D1
		inout  wire        hps_io_hps_io_usb1_inst_D2,                       //                       .hps_io_usb1_inst_D2
		inout  wire        hps_io_hps_io_usb1_inst_D3,                       //                       .hps_io_usb1_inst_D3
		inout  wire        hps_io_hps_io_usb1_inst_D4,                       //                       .hps_io_usb1_inst_D4
		inout  wire        hps_io_hps_io_usb1_inst_D5,                       //                       .hps_io_usb1_inst_D5
		inout  wire        hps_io_hps_io_usb1_inst_D6,                       //                       .hps_io_usb1_inst_D6
		inout  wire        hps_io_hps_io_usb1_inst_D7,                       //                       .hps_io_usb1_inst_D7
		input  wire        hps_io_hps_io_usb1_inst_CLK,                      //                       .hps_io_usb1_inst_CLK
		output wire        hps_io_hps_io_usb1_inst_STP,                      //                       .hps_io_usb1_inst_STP
		input  wire        hps_io_hps_io_usb1_inst_DIR,                      //                       .hps_io_usb1_inst_DIR
		input  wire        hps_io_hps_io_usb1_inst_NXT,                      //                       .hps_io_usb1_inst_NXT
		input  wire        hps_io_hps_io_uart0_inst_RX,                      //                       .hps_io_uart0_inst_RX
		output wire        hps_io_hps_io_uart0_inst_TX,                      //                       .hps_io_uart0_inst_TX
		inout  wire        hps_io_hps_io_i2c0_inst_SDA,                      //                       .hps_io_i2c0_inst_SDA
		inout  wire        hps_io_hps_io_i2c0_inst_SCL,                      //                       .hps_io_i2c0_inst_SCL
		inout  wire        hps_io_hps_io_gpio_inst_GPIO09,                   //                       .hps_io_gpio_inst_GPIO09
		inout  wire        hps_io_hps_io_gpio_inst_GPIO35,                   //                       .hps_io_gpio_inst_GPIO35
		inout  wire        hps_io_hps_io_gpio_inst_GPIO53,                   //                       .hps_io_gpio_inst_GPIO53
		inout  wire        hps_io_hps_io_gpio_inst_GPIO54,                   //                       .hps_io_gpio_inst_GPIO54
		inout  wire        hps_io_hps_io_gpio_inst_GPIO61,                   //                       .hps_io_gpio_inst_GPIO61
		output wire [14:0] hps_memory_mem_a,                                 //             hps_memory.mem_a
		output wire [2:0]  hps_memory_mem_ba,                                //                       .mem_ba
		output wire        hps_memory_mem_ck,                                //                       .mem_ck
		output wire        hps_memory_mem_ck_n,                              //                       .mem_ck_n
		output wire        hps_memory_mem_cke,                               //                       .mem_cke
		output wire        hps_memory_mem_cs_n,                              //                       .mem_cs_n
		output wire        hps_memory_mem_ras_n,                             //                       .mem_ras_n
		output wire        hps_memory_mem_cas_n,                             //                       .mem_cas_n
		output wire        hps_memory_mem_we_n,                              //                       .mem_we_n
		output wire        hps_memory_mem_reset_n,                           //                       .mem_reset_n
		inout  wire [31:0] hps_memory_mem_dq,                                //                       .mem_dq
		inout  wire [3:0]  hps_memory_mem_dqs,                               //                       .mem_dqs
		inout  wire [3:0]  hps_memory_mem_dqs_n,                             //                       .mem_dqs_n
		output wire        hps_memory_mem_odt,                               //                       .mem_odt
		output wire [3:0]  hps_memory_mem_dm,                                //                       .mem_dm
		input  wire        hps_memory_oct_rzqin,                             //                       .oct_rzqin
		input  wire        reset_reset_n                                     //                  reset.reset_n
	);

	wire   [1:0] hps_h2f_axi_master_awburst;                    // hps:h2f_AWBURST -> mm_interconnect_0:hps_h2f_axi_master_awburst
	wire   [3:0] hps_h2f_axi_master_arlen;                      // hps:h2f_ARLEN -> mm_interconnect_0:hps_h2f_axi_master_arlen
	wire   [3:0] hps_h2f_axi_master_wstrb;                      // hps:h2f_WSTRB -> mm_interconnect_0:hps_h2f_axi_master_wstrb
	wire         hps_h2f_axi_master_wready;                     // mm_interconnect_0:hps_h2f_axi_master_wready -> hps:h2f_WREADY
	wire  [11:0] hps_h2f_axi_master_rid;                        // mm_interconnect_0:hps_h2f_axi_master_rid -> hps:h2f_RID
	wire         hps_h2f_axi_master_rready;                     // hps:h2f_RREADY -> mm_interconnect_0:hps_h2f_axi_master_rready
	wire   [3:0] hps_h2f_axi_master_awlen;                      // hps:h2f_AWLEN -> mm_interconnect_0:hps_h2f_axi_master_awlen
	wire  [11:0] hps_h2f_axi_master_wid;                        // hps:h2f_WID -> mm_interconnect_0:hps_h2f_axi_master_wid
	wire   [3:0] hps_h2f_axi_master_arcache;                    // hps:h2f_ARCACHE -> mm_interconnect_0:hps_h2f_axi_master_arcache
	wire         hps_h2f_axi_master_wvalid;                     // hps:h2f_WVALID -> mm_interconnect_0:hps_h2f_axi_master_wvalid
	wire  [29:0] hps_h2f_axi_master_araddr;                     // hps:h2f_ARADDR -> mm_interconnect_0:hps_h2f_axi_master_araddr
	wire   [2:0] hps_h2f_axi_master_arprot;                     // hps:h2f_ARPROT -> mm_interconnect_0:hps_h2f_axi_master_arprot
	wire   [2:0] hps_h2f_axi_master_awprot;                     // hps:h2f_AWPROT -> mm_interconnect_0:hps_h2f_axi_master_awprot
	wire  [31:0] hps_h2f_axi_master_wdata;                      // hps:h2f_WDATA -> mm_interconnect_0:hps_h2f_axi_master_wdata
	wire         hps_h2f_axi_master_arvalid;                    // hps:h2f_ARVALID -> mm_interconnect_0:hps_h2f_axi_master_arvalid
	wire   [3:0] hps_h2f_axi_master_awcache;                    // hps:h2f_AWCACHE -> mm_interconnect_0:hps_h2f_axi_master_awcache
	wire  [11:0] hps_h2f_axi_master_arid;                       // hps:h2f_ARID -> mm_interconnect_0:hps_h2f_axi_master_arid
	wire   [1:0] hps_h2f_axi_master_arlock;                     // hps:h2f_ARLOCK -> mm_interconnect_0:hps_h2f_axi_master_arlock
	wire   [1:0] hps_h2f_axi_master_awlock;                     // hps:h2f_AWLOCK -> mm_interconnect_0:hps_h2f_axi_master_awlock
	wire  [29:0] hps_h2f_axi_master_awaddr;                     // hps:h2f_AWADDR -> mm_interconnect_0:hps_h2f_axi_master_awaddr
	wire   [1:0] hps_h2f_axi_master_bresp;                      // mm_interconnect_0:hps_h2f_axi_master_bresp -> hps:h2f_BRESP
	wire         hps_h2f_axi_master_arready;                    // mm_interconnect_0:hps_h2f_axi_master_arready -> hps:h2f_ARREADY
	wire  [31:0] hps_h2f_axi_master_rdata;                      // mm_interconnect_0:hps_h2f_axi_master_rdata -> hps:h2f_RDATA
	wire         hps_h2f_axi_master_awready;                    // mm_interconnect_0:hps_h2f_axi_master_awready -> hps:h2f_AWREADY
	wire   [1:0] hps_h2f_axi_master_arburst;                    // hps:h2f_ARBURST -> mm_interconnect_0:hps_h2f_axi_master_arburst
	wire   [2:0] hps_h2f_axi_master_arsize;                     // hps:h2f_ARSIZE -> mm_interconnect_0:hps_h2f_axi_master_arsize
	wire         hps_h2f_axi_master_bready;                     // hps:h2f_BREADY -> mm_interconnect_0:hps_h2f_axi_master_bready
	wire         hps_h2f_axi_master_rlast;                      // mm_interconnect_0:hps_h2f_axi_master_rlast -> hps:h2f_RLAST
	wire         hps_h2f_axi_master_wlast;                      // hps:h2f_WLAST -> mm_interconnect_0:hps_h2f_axi_master_wlast
	wire   [1:0] hps_h2f_axi_master_rresp;                      // mm_interconnect_0:hps_h2f_axi_master_rresp -> hps:h2f_RRESP
	wire  [11:0] hps_h2f_axi_master_awid;                       // hps:h2f_AWID -> mm_interconnect_0:hps_h2f_axi_master_awid
	wire  [11:0] hps_h2f_axi_master_bid;                        // mm_interconnect_0:hps_h2f_axi_master_bid -> hps:h2f_BID
	wire         hps_h2f_axi_master_bvalid;                     // mm_interconnect_0:hps_h2f_axi_master_bvalid -> hps:h2f_BVALID
	wire   [2:0] hps_h2f_axi_master_awsize;                     // hps:h2f_AWSIZE -> mm_interconnect_0:hps_h2f_axi_master_awsize
	wire         hps_h2f_axi_master_awvalid;                    // hps:h2f_AWVALID -> mm_interconnect_0:hps_h2f_axi_master_awvalid
	wire         hps_h2f_axi_master_rvalid;                     // mm_interconnect_0:hps_h2f_axi_master_rvalid -> hps:h2f_RVALID
	wire   [1:0] hps_h2f_lw_axi_master_awburst;                 // hps:h2f_lw_AWBURST -> mm_interconnect_0:hps_h2f_lw_axi_master_awburst
	wire   [3:0] hps_h2f_lw_axi_master_arlen;                   // hps:h2f_lw_ARLEN -> mm_interconnect_0:hps_h2f_lw_axi_master_arlen
	wire   [3:0] hps_h2f_lw_axi_master_wstrb;                   // hps:h2f_lw_WSTRB -> mm_interconnect_0:hps_h2f_lw_axi_master_wstrb
	wire         hps_h2f_lw_axi_master_wready;                  // mm_interconnect_0:hps_h2f_lw_axi_master_wready -> hps:h2f_lw_WREADY
	wire  [11:0] hps_h2f_lw_axi_master_rid;                     // mm_interconnect_0:hps_h2f_lw_axi_master_rid -> hps:h2f_lw_RID
	wire         hps_h2f_lw_axi_master_rready;                  // hps:h2f_lw_RREADY -> mm_interconnect_0:hps_h2f_lw_axi_master_rready
	wire   [3:0] hps_h2f_lw_axi_master_awlen;                   // hps:h2f_lw_AWLEN -> mm_interconnect_0:hps_h2f_lw_axi_master_awlen
	wire  [11:0] hps_h2f_lw_axi_master_wid;                     // hps:h2f_lw_WID -> mm_interconnect_0:hps_h2f_lw_axi_master_wid
	wire   [3:0] hps_h2f_lw_axi_master_arcache;                 // hps:h2f_lw_ARCACHE -> mm_interconnect_0:hps_h2f_lw_axi_master_arcache
	wire         hps_h2f_lw_axi_master_wvalid;                  // hps:h2f_lw_WVALID -> mm_interconnect_0:hps_h2f_lw_axi_master_wvalid
	wire  [20:0] hps_h2f_lw_axi_master_araddr;                  // hps:h2f_lw_ARADDR -> mm_interconnect_0:hps_h2f_lw_axi_master_araddr
	wire   [2:0] hps_h2f_lw_axi_master_arprot;                  // hps:h2f_lw_ARPROT -> mm_interconnect_0:hps_h2f_lw_axi_master_arprot
	wire   [2:0] hps_h2f_lw_axi_master_awprot;                  // hps:h2f_lw_AWPROT -> mm_interconnect_0:hps_h2f_lw_axi_master_awprot
	wire  [31:0] hps_h2f_lw_axi_master_wdata;                   // hps:h2f_lw_WDATA -> mm_interconnect_0:hps_h2f_lw_axi_master_wdata
	wire         hps_h2f_lw_axi_master_arvalid;                 // hps:h2f_lw_ARVALID -> mm_interconnect_0:hps_h2f_lw_axi_master_arvalid
	wire   [3:0] hps_h2f_lw_axi_master_awcache;                 // hps:h2f_lw_AWCACHE -> mm_interconnect_0:hps_h2f_lw_axi_master_awcache
	wire  [11:0] hps_h2f_lw_axi_master_arid;                    // hps:h2f_lw_ARID -> mm_interconnect_0:hps_h2f_lw_axi_master_arid
	wire   [1:0] hps_h2f_lw_axi_master_arlock;                  // hps:h2f_lw_ARLOCK -> mm_interconnect_0:hps_h2f_lw_axi_master_arlock
	wire   [1:0] hps_h2f_lw_axi_master_awlock;                  // hps:h2f_lw_AWLOCK -> mm_interconnect_0:hps_h2f_lw_axi_master_awlock
	wire  [20:0] hps_h2f_lw_axi_master_awaddr;                  // hps:h2f_lw_AWADDR -> mm_interconnect_0:hps_h2f_lw_axi_master_awaddr
	wire   [1:0] hps_h2f_lw_axi_master_bresp;                   // mm_interconnect_0:hps_h2f_lw_axi_master_bresp -> hps:h2f_lw_BRESP
	wire         hps_h2f_lw_axi_master_arready;                 // mm_interconnect_0:hps_h2f_lw_axi_master_arready -> hps:h2f_lw_ARREADY
	wire  [31:0] hps_h2f_lw_axi_master_rdata;                   // mm_interconnect_0:hps_h2f_lw_axi_master_rdata -> hps:h2f_lw_RDATA
	wire         hps_h2f_lw_axi_master_awready;                 // mm_interconnect_0:hps_h2f_lw_axi_master_awready -> hps:h2f_lw_AWREADY
	wire   [1:0] hps_h2f_lw_axi_master_arburst;                 // hps:h2f_lw_ARBURST -> mm_interconnect_0:hps_h2f_lw_axi_master_arburst
	wire   [2:0] hps_h2f_lw_axi_master_arsize;                  // hps:h2f_lw_ARSIZE -> mm_interconnect_0:hps_h2f_lw_axi_master_arsize
	wire         hps_h2f_lw_axi_master_bready;                  // hps:h2f_lw_BREADY -> mm_interconnect_0:hps_h2f_lw_axi_master_bready
	wire         hps_h2f_lw_axi_master_rlast;                   // mm_interconnect_0:hps_h2f_lw_axi_master_rlast -> hps:h2f_lw_RLAST
	wire         hps_h2f_lw_axi_master_wlast;                   // hps:h2f_lw_WLAST -> mm_interconnect_0:hps_h2f_lw_axi_master_wlast
	wire   [1:0] hps_h2f_lw_axi_master_rresp;                   // mm_interconnect_0:hps_h2f_lw_axi_master_rresp -> hps:h2f_lw_RRESP
	wire  [11:0] hps_h2f_lw_axi_master_awid;                    // hps:h2f_lw_AWID -> mm_interconnect_0:hps_h2f_lw_axi_master_awid
	wire  [11:0] hps_h2f_lw_axi_master_bid;                     // mm_interconnect_0:hps_h2f_lw_axi_master_bid -> hps:h2f_lw_BID
	wire         hps_h2f_lw_axi_master_bvalid;                  // mm_interconnect_0:hps_h2f_lw_axi_master_bvalid -> hps:h2f_lw_BVALID
	wire   [2:0] hps_h2f_lw_axi_master_awsize;                  // hps:h2f_lw_AWSIZE -> mm_interconnect_0:hps_h2f_lw_axi_master_awsize
	wire         hps_h2f_lw_axi_master_awvalid;                 // hps:h2f_lw_AWVALID -> mm_interconnect_0:hps_h2f_lw_axi_master_awvalid
	wire         hps_h2f_lw_axi_master_rvalid;                  // mm_interconnect_0:hps_h2f_lw_axi_master_rvalid -> hps:h2f_lw_RVALID
	wire         mm_interconnect_0_onchip_memory_s1_chipselect; // mm_interconnect_0:onchip_memory_s1_chipselect -> onchip_memory:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_readdata;   // onchip_memory:readdata -> mm_interconnect_0:onchip_memory_s1_readdata
	wire  [11:0] mm_interconnect_0_onchip_memory_s1_address;    // mm_interconnect_0:onchip_memory_s1_address -> onchip_memory:address
	wire   [3:0] mm_interconnect_0_onchip_memory_s1_byteenable; // mm_interconnect_0:onchip_memory_s1_byteenable -> onchip_memory:byteenable
	wire         mm_interconnect_0_onchip_memory_s1_write;      // mm_interconnect_0:onchip_memory_s1_write -> onchip_memory:write
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_writedata;  // mm_interconnect_0:onchip_memory_s1_writedata -> onchip_memory:writedata
	wire         mm_interconnect_0_onchip_memory_s1_clken;      // mm_interconnect_0:onchip_memory_s1_clken -> onchip_memory:clken
	wire  [31:0] hps_f2h_irq0_irq;                              // irq_mapper:sender_irq -> hps:f2h_irq_p0
	wire  [31:0] hps_f2h_irq1_irq;                              // irq_mapper_001:sender_irq -> hps:f2h_irq_p1
	wire         rst_controller_reset_out_reset;                // rst_controller:reset_out -> [mm_interconnect_0:onchip_memory_reset1_reset_bridge_in_reset_reset, onchip_memory:reset]
	wire         rst_controller_001_reset_out_reset;            // rst_controller_001:reset_out -> mm_interconnect_0:hps_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset

	HPS_hps #(
		.F2S_Width (1),
		.S2F_Width (1)
	) hps (
		.f2h_boot_from_fpga_ready      (hps_f2h_boot_from_fpga_boot_from_fpga_ready),      // f2h_boot_from_fpga.boot_from_fpga_ready
		.f2h_boot_from_fpga_on_failure (hps_f2h_boot_from_fpga_boot_from_fpga_on_failure), //                   .boot_from_fpga_on_failure
		.mem_a                         (hps_memory_mem_a),                                 //             memory.mem_a
		.mem_ba                        (hps_memory_mem_ba),                                //                   .mem_ba
		.mem_ck                        (hps_memory_mem_ck),                                //                   .mem_ck
		.mem_ck_n                      (hps_memory_mem_ck_n),                              //                   .mem_ck_n
		.mem_cke                       (hps_memory_mem_cke),                               //                   .mem_cke
		.mem_cs_n                      (hps_memory_mem_cs_n),                              //                   .mem_cs_n
		.mem_ras_n                     (hps_memory_mem_ras_n),                             //                   .mem_ras_n
		.mem_cas_n                     (hps_memory_mem_cas_n),                             //                   .mem_cas_n
		.mem_we_n                      (hps_memory_mem_we_n),                              //                   .mem_we_n
		.mem_reset_n                   (hps_memory_mem_reset_n),                           //                   .mem_reset_n
		.mem_dq                        (hps_memory_mem_dq),                                //                   .mem_dq
		.mem_dqs                       (hps_memory_mem_dqs),                               //                   .mem_dqs
		.mem_dqs_n                     (hps_memory_mem_dqs_n),                             //                   .mem_dqs_n
		.mem_odt                       (hps_memory_mem_odt),                               //                   .mem_odt
		.mem_dm                        (hps_memory_mem_dm),                                //                   .mem_dm
		.oct_rzqin                     (hps_memory_oct_rzqin),                             //                   .oct_rzqin
		.hps_io_emac1_inst_TX_CLK      (hps_io_hps_io_emac1_inst_TX_CLK),                  //             hps_io.hps_io_emac1_inst_TX_CLK
		.hps_io_emac1_inst_TXD0        (hps_io_hps_io_emac1_inst_TXD0),                    //                   .hps_io_emac1_inst_TXD0
		.hps_io_emac1_inst_TXD1        (hps_io_hps_io_emac1_inst_TXD1),                    //                   .hps_io_emac1_inst_TXD1
		.hps_io_emac1_inst_TXD2        (hps_io_hps_io_emac1_inst_TXD2),                    //                   .hps_io_emac1_inst_TXD2
		.hps_io_emac1_inst_TXD3        (hps_io_hps_io_emac1_inst_TXD3),                    //                   .hps_io_emac1_inst_TXD3
		.hps_io_emac1_inst_RXD0        (hps_io_hps_io_emac1_inst_RXD0),                    //                   .hps_io_emac1_inst_RXD0
		.hps_io_emac1_inst_MDIO        (hps_io_hps_io_emac1_inst_MDIO),                    //                   .hps_io_emac1_inst_MDIO
		.hps_io_emac1_inst_MDC         (hps_io_hps_io_emac1_inst_MDC),                     //                   .hps_io_emac1_inst_MDC
		.hps_io_emac1_inst_RX_CTL      (hps_io_hps_io_emac1_inst_RX_CTL),                  //                   .hps_io_emac1_inst_RX_CTL
		.hps_io_emac1_inst_TX_CTL      (hps_io_hps_io_emac1_inst_TX_CTL),                  //                   .hps_io_emac1_inst_TX_CTL
		.hps_io_emac1_inst_RX_CLK      (hps_io_hps_io_emac1_inst_RX_CLK),                  //                   .hps_io_emac1_inst_RX_CLK
		.hps_io_emac1_inst_RXD1        (hps_io_hps_io_emac1_inst_RXD1),                    //                   .hps_io_emac1_inst_RXD1
		.hps_io_emac1_inst_RXD2        (hps_io_hps_io_emac1_inst_RXD2),                    //                   .hps_io_emac1_inst_RXD2
		.hps_io_emac1_inst_RXD3        (hps_io_hps_io_emac1_inst_RXD3),                    //                   .hps_io_emac1_inst_RXD3
		.hps_io_sdio_inst_CMD          (hps_io_hps_io_sdio_inst_CMD),                      //                   .hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0           (hps_io_hps_io_sdio_inst_D0),                       //                   .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1           (hps_io_hps_io_sdio_inst_D1),                       //                   .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_CLK          (hps_io_hps_io_sdio_inst_CLK),                      //                   .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2           (hps_io_hps_io_sdio_inst_D2),                       //                   .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3           (hps_io_hps_io_sdio_inst_D3),                       //                   .hps_io_sdio_inst_D3
		.hps_io_usb1_inst_D0           (hps_io_hps_io_usb1_inst_D0),                       //                   .hps_io_usb1_inst_D0
		.hps_io_usb1_inst_D1           (hps_io_hps_io_usb1_inst_D1),                       //                   .hps_io_usb1_inst_D1
		.hps_io_usb1_inst_D2           (hps_io_hps_io_usb1_inst_D2),                       //                   .hps_io_usb1_inst_D2
		.hps_io_usb1_inst_D3           (hps_io_hps_io_usb1_inst_D3),                       //                   .hps_io_usb1_inst_D3
		.hps_io_usb1_inst_D4           (hps_io_hps_io_usb1_inst_D4),                       //                   .hps_io_usb1_inst_D4
		.hps_io_usb1_inst_D5           (hps_io_hps_io_usb1_inst_D5),                       //                   .hps_io_usb1_inst_D5
		.hps_io_usb1_inst_D6           (hps_io_hps_io_usb1_inst_D6),                       //                   .hps_io_usb1_inst_D6
		.hps_io_usb1_inst_D7           (hps_io_hps_io_usb1_inst_D7),                       //                   .hps_io_usb1_inst_D7
		.hps_io_usb1_inst_CLK          (hps_io_hps_io_usb1_inst_CLK),                      //                   .hps_io_usb1_inst_CLK
		.hps_io_usb1_inst_STP          (hps_io_hps_io_usb1_inst_STP),                      //                   .hps_io_usb1_inst_STP
		.hps_io_usb1_inst_DIR          (hps_io_hps_io_usb1_inst_DIR),                      //                   .hps_io_usb1_inst_DIR
		.hps_io_usb1_inst_NXT          (hps_io_hps_io_usb1_inst_NXT),                      //                   .hps_io_usb1_inst_NXT
		.hps_io_uart0_inst_RX          (hps_io_hps_io_uart0_inst_RX),                      //                   .hps_io_uart0_inst_RX
		.hps_io_uart0_inst_TX          (hps_io_hps_io_uart0_inst_TX),                      //                   .hps_io_uart0_inst_TX
		.hps_io_i2c0_inst_SDA          (hps_io_hps_io_i2c0_inst_SDA),                      //                   .hps_io_i2c0_inst_SDA
		.hps_io_i2c0_inst_SCL          (hps_io_hps_io_i2c0_inst_SCL),                      //                   .hps_io_i2c0_inst_SCL
		.hps_io_gpio_inst_GPIO09       (hps_io_hps_io_gpio_inst_GPIO09),                   //                   .hps_io_gpio_inst_GPIO09
		.hps_io_gpio_inst_GPIO35       (hps_io_hps_io_gpio_inst_GPIO35),                   //                   .hps_io_gpio_inst_GPIO35
		.hps_io_gpio_inst_GPIO53       (hps_io_hps_io_gpio_inst_GPIO53),                   //                   .hps_io_gpio_inst_GPIO53
		.hps_io_gpio_inst_GPIO54       (hps_io_hps_io_gpio_inst_GPIO54),                   //                   .hps_io_gpio_inst_GPIO54
		.hps_io_gpio_inst_GPIO61       (hps_io_hps_io_gpio_inst_GPIO61),                   //                   .hps_io_gpio_inst_GPIO61
		.h2f_rst_n                     (hps_h2f_reset_reset_n),                            //          h2f_reset.reset_n
		.h2f_axi_clk                   (clk_clk),                                          //      h2f_axi_clock.clk
		.h2f_AWID                      (hps_h2f_axi_master_awid),                          //     h2f_axi_master.awid
		.h2f_AWADDR                    (hps_h2f_axi_master_awaddr),                        //                   .awaddr
		.h2f_AWLEN                     (hps_h2f_axi_master_awlen),                         //                   .awlen
		.h2f_AWSIZE                    (hps_h2f_axi_master_awsize),                        //                   .awsize
		.h2f_AWBURST                   (hps_h2f_axi_master_awburst),                       //                   .awburst
		.h2f_AWLOCK                    (hps_h2f_axi_master_awlock),                        //                   .awlock
		.h2f_AWCACHE                   (hps_h2f_axi_master_awcache),                       //                   .awcache
		.h2f_AWPROT                    (hps_h2f_axi_master_awprot),                        //                   .awprot
		.h2f_AWVALID                   (hps_h2f_axi_master_awvalid),                       //                   .awvalid
		.h2f_AWREADY                   (hps_h2f_axi_master_awready),                       //                   .awready
		.h2f_WID                       (hps_h2f_axi_master_wid),                           //                   .wid
		.h2f_WDATA                     (hps_h2f_axi_master_wdata),                         //                   .wdata
		.h2f_WSTRB                     (hps_h2f_axi_master_wstrb),                         //                   .wstrb
		.h2f_WLAST                     (hps_h2f_axi_master_wlast),                         //                   .wlast
		.h2f_WVALID                    (hps_h2f_axi_master_wvalid),                        //                   .wvalid
		.h2f_WREADY                    (hps_h2f_axi_master_wready),                        //                   .wready
		.h2f_BID                       (hps_h2f_axi_master_bid),                           //                   .bid
		.h2f_BRESP                     (hps_h2f_axi_master_bresp),                         //                   .bresp
		.h2f_BVALID                    (hps_h2f_axi_master_bvalid),                        //                   .bvalid
		.h2f_BREADY                    (hps_h2f_axi_master_bready),                        //                   .bready
		.h2f_ARID                      (hps_h2f_axi_master_arid),                          //                   .arid
		.h2f_ARADDR                    (hps_h2f_axi_master_araddr),                        //                   .araddr
		.h2f_ARLEN                     (hps_h2f_axi_master_arlen),                         //                   .arlen
		.h2f_ARSIZE                    (hps_h2f_axi_master_arsize),                        //                   .arsize
		.h2f_ARBURST                   (hps_h2f_axi_master_arburst),                       //                   .arburst
		.h2f_ARLOCK                    (hps_h2f_axi_master_arlock),                        //                   .arlock
		.h2f_ARCACHE                   (hps_h2f_axi_master_arcache),                       //                   .arcache
		.h2f_ARPROT                    (hps_h2f_axi_master_arprot),                        //                   .arprot
		.h2f_ARVALID                   (hps_h2f_axi_master_arvalid),                       //                   .arvalid
		.h2f_ARREADY                   (hps_h2f_axi_master_arready),                       //                   .arready
		.h2f_RID                       (hps_h2f_axi_master_rid),                           //                   .rid
		.h2f_RDATA                     (hps_h2f_axi_master_rdata),                         //                   .rdata
		.h2f_RRESP                     (hps_h2f_axi_master_rresp),                         //                   .rresp
		.h2f_RLAST                     (hps_h2f_axi_master_rlast),                         //                   .rlast
		.h2f_RVALID                    (hps_h2f_axi_master_rvalid),                        //                   .rvalid
		.h2f_RREADY                    (hps_h2f_axi_master_rready),                        //                   .rready
		.f2h_axi_clk                   (hps_f2h_axi_clock_clk),                            //      f2h_axi_clock.clk
		.f2h_AWID                      (hps_f2h_axi_slave_awid),                           //      f2h_axi_slave.awid
		.f2h_AWADDR                    (hps_f2h_axi_slave_awaddr),                         //                   .awaddr
		.f2h_AWLEN                     (hps_f2h_axi_slave_awlen),                          //                   .awlen
		.f2h_AWSIZE                    (hps_f2h_axi_slave_awsize),                         //                   .awsize
		.f2h_AWBURST                   (hps_f2h_axi_slave_awburst),                        //                   .awburst
		.f2h_AWLOCK                    (hps_f2h_axi_slave_awlock),                         //                   .awlock
		.f2h_AWCACHE                   (hps_f2h_axi_slave_awcache),                        //                   .awcache
		.f2h_AWPROT                    (hps_f2h_axi_slave_awprot),                         //                   .awprot
		.f2h_AWVALID                   (hps_f2h_axi_slave_awvalid),                        //                   .awvalid
		.f2h_AWREADY                   (hps_f2h_axi_slave_awready),                        //                   .awready
		.f2h_AWUSER                    (hps_f2h_axi_slave_awuser),                         //                   .awuser
		.f2h_WID                       (hps_f2h_axi_slave_wid),                            //                   .wid
		.f2h_WDATA                     (hps_f2h_axi_slave_wdata),                          //                   .wdata
		.f2h_WSTRB                     (hps_f2h_axi_slave_wstrb),                          //                   .wstrb
		.f2h_WLAST                     (hps_f2h_axi_slave_wlast),                          //                   .wlast
		.f2h_WVALID                    (hps_f2h_axi_slave_wvalid),                         //                   .wvalid
		.f2h_WREADY                    (hps_f2h_axi_slave_wready),                         //                   .wready
		.f2h_BID                       (hps_f2h_axi_slave_bid),                            //                   .bid
		.f2h_BRESP                     (hps_f2h_axi_slave_bresp),                          //                   .bresp
		.f2h_BVALID                    (hps_f2h_axi_slave_bvalid),                         //                   .bvalid
		.f2h_BREADY                    (hps_f2h_axi_slave_bready),                         //                   .bready
		.f2h_ARID                      (hps_f2h_axi_slave_arid),                           //                   .arid
		.f2h_ARADDR                    (hps_f2h_axi_slave_araddr),                         //                   .araddr
		.f2h_ARLEN                     (hps_f2h_axi_slave_arlen),                          //                   .arlen
		.f2h_ARSIZE                    (hps_f2h_axi_slave_arsize),                         //                   .arsize
		.f2h_ARBURST                   (hps_f2h_axi_slave_arburst),                        //                   .arburst
		.f2h_ARLOCK                    (hps_f2h_axi_slave_arlock),                         //                   .arlock
		.f2h_ARCACHE                   (hps_f2h_axi_slave_arcache),                        //                   .arcache
		.f2h_ARPROT                    (hps_f2h_axi_slave_arprot),                         //                   .arprot
		.f2h_ARVALID                   (hps_f2h_axi_slave_arvalid),                        //                   .arvalid
		.f2h_ARREADY                   (hps_f2h_axi_slave_arready),                        //                   .arready
		.f2h_ARUSER                    (hps_f2h_axi_slave_aruser),                         //                   .aruser
		.f2h_RID                       (hps_f2h_axi_slave_rid),                            //                   .rid
		.f2h_RDATA                     (hps_f2h_axi_slave_rdata),                          //                   .rdata
		.f2h_RRESP                     (hps_f2h_axi_slave_rresp),                          //                   .rresp
		.f2h_RLAST                     (hps_f2h_axi_slave_rlast),                          //                   .rlast
		.f2h_RVALID                    (hps_f2h_axi_slave_rvalid),                         //                   .rvalid
		.f2h_RREADY                    (hps_f2h_axi_slave_rready),                         //                   .rready
		.h2f_lw_axi_clk                (clk_clk),                                          //   h2f_lw_axi_clock.clk
		.h2f_lw_AWID                   (hps_h2f_lw_axi_master_awid),                       //  h2f_lw_axi_master.awid
		.h2f_lw_AWADDR                 (hps_h2f_lw_axi_master_awaddr),                     //                   .awaddr
		.h2f_lw_AWLEN                  (hps_h2f_lw_axi_master_awlen),                      //                   .awlen
		.h2f_lw_AWSIZE                 (hps_h2f_lw_axi_master_awsize),                     //                   .awsize
		.h2f_lw_AWBURST                (hps_h2f_lw_axi_master_awburst),                    //                   .awburst
		.h2f_lw_AWLOCK                 (hps_h2f_lw_axi_master_awlock),                     //                   .awlock
		.h2f_lw_AWCACHE                (hps_h2f_lw_axi_master_awcache),                    //                   .awcache
		.h2f_lw_AWPROT                 (hps_h2f_lw_axi_master_awprot),                     //                   .awprot
		.h2f_lw_AWVALID                (hps_h2f_lw_axi_master_awvalid),                    //                   .awvalid
		.h2f_lw_AWREADY                (hps_h2f_lw_axi_master_awready),                    //                   .awready
		.h2f_lw_WID                    (hps_h2f_lw_axi_master_wid),                        //                   .wid
		.h2f_lw_WDATA                  (hps_h2f_lw_axi_master_wdata),                      //                   .wdata
		.h2f_lw_WSTRB                  (hps_h2f_lw_axi_master_wstrb),                      //                   .wstrb
		.h2f_lw_WLAST                  (hps_h2f_lw_axi_master_wlast),                      //                   .wlast
		.h2f_lw_WVALID                 (hps_h2f_lw_axi_master_wvalid),                     //                   .wvalid
		.h2f_lw_WREADY                 (hps_h2f_lw_axi_master_wready),                     //                   .wready
		.h2f_lw_BID                    (hps_h2f_lw_axi_master_bid),                        //                   .bid
		.h2f_lw_BRESP                  (hps_h2f_lw_axi_master_bresp),                      //                   .bresp
		.h2f_lw_BVALID                 (hps_h2f_lw_axi_master_bvalid),                     //                   .bvalid
		.h2f_lw_BREADY                 (hps_h2f_lw_axi_master_bready),                     //                   .bready
		.h2f_lw_ARID                   (hps_h2f_lw_axi_master_arid),                       //                   .arid
		.h2f_lw_ARADDR                 (hps_h2f_lw_axi_master_araddr),                     //                   .araddr
		.h2f_lw_ARLEN                  (hps_h2f_lw_axi_master_arlen),                      //                   .arlen
		.h2f_lw_ARSIZE                 (hps_h2f_lw_axi_master_arsize),                     //                   .arsize
		.h2f_lw_ARBURST                (hps_h2f_lw_axi_master_arburst),                    //                   .arburst
		.h2f_lw_ARLOCK                 (hps_h2f_lw_axi_master_arlock),                     //                   .arlock
		.h2f_lw_ARCACHE                (hps_h2f_lw_axi_master_arcache),                    //                   .arcache
		.h2f_lw_ARPROT                 (hps_h2f_lw_axi_master_arprot),                     //                   .arprot
		.h2f_lw_ARVALID                (hps_h2f_lw_axi_master_arvalid),                    //                   .arvalid
		.h2f_lw_ARREADY                (hps_h2f_lw_axi_master_arready),                    //                   .arready
		.h2f_lw_RID                    (hps_h2f_lw_axi_master_rid),                        //                   .rid
		.h2f_lw_RDATA                  (hps_h2f_lw_axi_master_rdata),                      //                   .rdata
		.h2f_lw_RRESP                  (hps_h2f_lw_axi_master_rresp),                      //                   .rresp
		.h2f_lw_RLAST                  (hps_h2f_lw_axi_master_rlast),                      //                   .rlast
		.h2f_lw_RVALID                 (hps_h2f_lw_axi_master_rvalid),                     //                   .rvalid
		.h2f_lw_RREADY                 (hps_h2f_lw_axi_master_rready),                     //                   .rready
		.f2h_irq_p0                    (hps_f2h_irq0_irq),                                 //           f2h_irq0.irq
		.f2h_irq_p1                    (hps_f2h_irq1_irq)                                  //           f2h_irq1.irq
	);

	HPS_onchip_memory onchip_memory (
		.clk        (clk_clk),                                       //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                // reset1.reset
		.reset_req  (1'b0),                                          // (terminated)
		.freeze     (1'b0)                                           // (terminated)
	);

	HPS_mm_interconnect_0 mm_interconnect_0 (
		.hps_h2f_axi_master_awid                                        (hps_h2f_axi_master_awid),                       //                                       hps_h2f_axi_master.awid
		.hps_h2f_axi_master_awaddr                                      (hps_h2f_axi_master_awaddr),                     //                                                         .awaddr
		.hps_h2f_axi_master_awlen                                       (hps_h2f_axi_master_awlen),                      //                                                         .awlen
		.hps_h2f_axi_master_awsize                                      (hps_h2f_axi_master_awsize),                     //                                                         .awsize
		.hps_h2f_axi_master_awburst                                     (hps_h2f_axi_master_awburst),                    //                                                         .awburst
		.hps_h2f_axi_master_awlock                                      (hps_h2f_axi_master_awlock),                     //                                                         .awlock
		.hps_h2f_axi_master_awcache                                     (hps_h2f_axi_master_awcache),                    //                                                         .awcache
		.hps_h2f_axi_master_awprot                                      (hps_h2f_axi_master_awprot),                     //                                                         .awprot
		.hps_h2f_axi_master_awvalid                                     (hps_h2f_axi_master_awvalid),                    //                                                         .awvalid
		.hps_h2f_axi_master_awready                                     (hps_h2f_axi_master_awready),                    //                                                         .awready
		.hps_h2f_axi_master_wid                                         (hps_h2f_axi_master_wid),                        //                                                         .wid
		.hps_h2f_axi_master_wdata                                       (hps_h2f_axi_master_wdata),                      //                                                         .wdata
		.hps_h2f_axi_master_wstrb                                       (hps_h2f_axi_master_wstrb),                      //                                                         .wstrb
		.hps_h2f_axi_master_wlast                                       (hps_h2f_axi_master_wlast),                      //                                                         .wlast
		.hps_h2f_axi_master_wvalid                                      (hps_h2f_axi_master_wvalid),                     //                                                         .wvalid
		.hps_h2f_axi_master_wready                                      (hps_h2f_axi_master_wready),                     //                                                         .wready
		.hps_h2f_axi_master_bid                                         (hps_h2f_axi_master_bid),                        //                                                         .bid
		.hps_h2f_axi_master_bresp                                       (hps_h2f_axi_master_bresp),                      //                                                         .bresp
		.hps_h2f_axi_master_bvalid                                      (hps_h2f_axi_master_bvalid),                     //                                                         .bvalid
		.hps_h2f_axi_master_bready                                      (hps_h2f_axi_master_bready),                     //                                                         .bready
		.hps_h2f_axi_master_arid                                        (hps_h2f_axi_master_arid),                       //                                                         .arid
		.hps_h2f_axi_master_araddr                                      (hps_h2f_axi_master_araddr),                     //                                                         .araddr
		.hps_h2f_axi_master_arlen                                       (hps_h2f_axi_master_arlen),                      //                                                         .arlen
		.hps_h2f_axi_master_arsize                                      (hps_h2f_axi_master_arsize),                     //                                                         .arsize
		.hps_h2f_axi_master_arburst                                     (hps_h2f_axi_master_arburst),                    //                                                         .arburst
		.hps_h2f_axi_master_arlock                                      (hps_h2f_axi_master_arlock),                     //                                                         .arlock
		.hps_h2f_axi_master_arcache                                     (hps_h2f_axi_master_arcache),                    //                                                         .arcache
		.hps_h2f_axi_master_arprot                                      (hps_h2f_axi_master_arprot),                     //                                                         .arprot
		.hps_h2f_axi_master_arvalid                                     (hps_h2f_axi_master_arvalid),                    //                                                         .arvalid
		.hps_h2f_axi_master_arready                                     (hps_h2f_axi_master_arready),                    //                                                         .arready
		.hps_h2f_axi_master_rid                                         (hps_h2f_axi_master_rid),                        //                                                         .rid
		.hps_h2f_axi_master_rdata                                       (hps_h2f_axi_master_rdata),                      //                                                         .rdata
		.hps_h2f_axi_master_rresp                                       (hps_h2f_axi_master_rresp),                      //                                                         .rresp
		.hps_h2f_axi_master_rlast                                       (hps_h2f_axi_master_rlast),                      //                                                         .rlast
		.hps_h2f_axi_master_rvalid                                      (hps_h2f_axi_master_rvalid),                     //                                                         .rvalid
		.hps_h2f_axi_master_rready                                      (hps_h2f_axi_master_rready),                     //                                                         .rready
		.hps_h2f_lw_axi_master_awid                                     (hps_h2f_lw_axi_master_awid),                    //                                    hps_h2f_lw_axi_master.awid
		.hps_h2f_lw_axi_master_awaddr                                   (hps_h2f_lw_axi_master_awaddr),                  //                                                         .awaddr
		.hps_h2f_lw_axi_master_awlen                                    (hps_h2f_lw_axi_master_awlen),                   //                                                         .awlen
		.hps_h2f_lw_axi_master_awsize                                   (hps_h2f_lw_axi_master_awsize),                  //                                                         .awsize
		.hps_h2f_lw_axi_master_awburst                                  (hps_h2f_lw_axi_master_awburst),                 //                                                         .awburst
		.hps_h2f_lw_axi_master_awlock                                   (hps_h2f_lw_axi_master_awlock),                  //                                                         .awlock
		.hps_h2f_lw_axi_master_awcache                                  (hps_h2f_lw_axi_master_awcache),                 //                                                         .awcache
		.hps_h2f_lw_axi_master_awprot                                   (hps_h2f_lw_axi_master_awprot),                  //                                                         .awprot
		.hps_h2f_lw_axi_master_awvalid                                  (hps_h2f_lw_axi_master_awvalid),                 //                                                         .awvalid
		.hps_h2f_lw_axi_master_awready                                  (hps_h2f_lw_axi_master_awready),                 //                                                         .awready
		.hps_h2f_lw_axi_master_wid                                      (hps_h2f_lw_axi_master_wid),                     //                                                         .wid
		.hps_h2f_lw_axi_master_wdata                                    (hps_h2f_lw_axi_master_wdata),                   //                                                         .wdata
		.hps_h2f_lw_axi_master_wstrb                                    (hps_h2f_lw_axi_master_wstrb),                   //                                                         .wstrb
		.hps_h2f_lw_axi_master_wlast                                    (hps_h2f_lw_axi_master_wlast),                   //                                                         .wlast
		.hps_h2f_lw_axi_master_wvalid                                   (hps_h2f_lw_axi_master_wvalid),                  //                                                         .wvalid
		.hps_h2f_lw_axi_master_wready                                   (hps_h2f_lw_axi_master_wready),                  //                                                         .wready
		.hps_h2f_lw_axi_master_bid                                      (hps_h2f_lw_axi_master_bid),                     //                                                         .bid
		.hps_h2f_lw_axi_master_bresp                                    (hps_h2f_lw_axi_master_bresp),                   //                                                         .bresp
		.hps_h2f_lw_axi_master_bvalid                                   (hps_h2f_lw_axi_master_bvalid),                  //                                                         .bvalid
		.hps_h2f_lw_axi_master_bready                                   (hps_h2f_lw_axi_master_bready),                  //                                                         .bready
		.hps_h2f_lw_axi_master_arid                                     (hps_h2f_lw_axi_master_arid),                    //                                                         .arid
		.hps_h2f_lw_axi_master_araddr                                   (hps_h2f_lw_axi_master_araddr),                  //                                                         .araddr
		.hps_h2f_lw_axi_master_arlen                                    (hps_h2f_lw_axi_master_arlen),                   //                                                         .arlen
		.hps_h2f_lw_axi_master_arsize                                   (hps_h2f_lw_axi_master_arsize),                  //                                                         .arsize
		.hps_h2f_lw_axi_master_arburst                                  (hps_h2f_lw_axi_master_arburst),                 //                                                         .arburst
		.hps_h2f_lw_axi_master_arlock                                   (hps_h2f_lw_axi_master_arlock),                  //                                                         .arlock
		.hps_h2f_lw_axi_master_arcache                                  (hps_h2f_lw_axi_master_arcache),                 //                                                         .arcache
		.hps_h2f_lw_axi_master_arprot                                   (hps_h2f_lw_axi_master_arprot),                  //                                                         .arprot
		.hps_h2f_lw_axi_master_arvalid                                  (hps_h2f_lw_axi_master_arvalid),                 //                                                         .arvalid
		.hps_h2f_lw_axi_master_arready                                  (hps_h2f_lw_axi_master_arready),                 //                                                         .arready
		.hps_h2f_lw_axi_master_rid                                      (hps_h2f_lw_axi_master_rid),                     //                                                         .rid
		.hps_h2f_lw_axi_master_rdata                                    (hps_h2f_lw_axi_master_rdata),                   //                                                         .rdata
		.hps_h2f_lw_axi_master_rresp                                    (hps_h2f_lw_axi_master_rresp),                   //                                                         .rresp
		.hps_h2f_lw_axi_master_rlast                                    (hps_h2f_lw_axi_master_rlast),                   //                                                         .rlast
		.hps_h2f_lw_axi_master_rvalid                                   (hps_h2f_lw_axi_master_rvalid),                  //                                                         .rvalid
		.hps_h2f_lw_axi_master_rready                                   (hps_h2f_lw_axi_master_rready),                  //                                                         .rready
		.clk_clk_clk                                                    (clk_clk),                                       //                                                  clk_clk.clk
		.hps_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),            // hps_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.onchip_memory_reset1_reset_bridge_in_reset_reset               (rst_controller_reset_out_reset),                //               onchip_memory_reset1_reset_bridge_in_reset.reset
		.onchip_memory_s1_address                                       (mm_interconnect_0_onchip_memory_s1_address),    //                                         onchip_memory_s1.address
		.onchip_memory_s1_write                                         (mm_interconnect_0_onchip_memory_s1_write),      //                                                         .write
		.onchip_memory_s1_readdata                                      (mm_interconnect_0_onchip_memory_s1_readdata),   //                                                         .readdata
		.onchip_memory_s1_writedata                                     (mm_interconnect_0_onchip_memory_s1_writedata),  //                                                         .writedata
		.onchip_memory_s1_byteenable                                    (mm_interconnect_0_onchip_memory_s1_byteenable), //                                                         .byteenable
		.onchip_memory_s1_chipselect                                    (mm_interconnect_0_onchip_memory_s1_chipselect), //                                                         .chipselect
		.onchip_memory_s1_clken                                         (mm_interconnect_0_onchip_memory_s1_clken)       //                                                         .clken
	);

	HPS_irq_mapper irq_mapper (
		.clk        (),                 //       clk.clk
		.reset      (),                 // clk_reset.reset
		.sender_irq (hps_f2h_irq0_irq)  //    sender.irq
	);

	HPS_irq_mapper irq_mapper_001 (
		.clk        (),                 //       clk.clk
		.reset      (),                 // clk_reset.reset
		.sender_irq (hps_f2h_irq1_irq)  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~hps_h2f_reset_reset_n),             // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
